module and_gate (y_out,a_in,b_in);

input a_in , b_in;
output y_out;

and dut(y_out,a_in,b_in);

endmodule

